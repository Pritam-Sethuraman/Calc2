library verilog;
use verilog.vl_types.all;
entity calc2_test is
end calc2_test;
